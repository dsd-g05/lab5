-- Descp.
--
-- entity name: g05_lab5
--
-- Version 1.0
-- Author: Felix Dube; felix.dube@mail.mcgill.ca & Auguste Lalande; auguste.lalande@mail.mcgill.ca
-- Date: November 26, 2015

library ieee;
use ieee.std_logic_1164.all;

entity g05_lab5 is
	port (
        START, READY : in std_logic;
        MODE : in std_logic;
        CLK : in std_logic;
	);
end g05_lab5;

architecture behavior of g05_lab5 is


end behavior;